package save_state_consts;
    parameter int SSIDX_GLOBAL = 0;
    parameter int SSIDX_SCN_RAM_0_LO = 1;
    parameter int SSIDX_SCN_RAM_0_UP = 2;
    parameter int SSIDX_PRI_RAM_L = 3;
    parameter int SSIDX_PRI_RAM_H = 4;
    parameter int SSIDX_CPU_RAM = 5;
    parameter int SSIDX_SCN_0 = 6;
endpackage


