module TC0360PRI #(parameter SS_IDX=-1) (
    input clk,
    input ce_pixel,
    input reset,

    // CPU Interface
    input [15:0] cpu_din,
    output reg [15:0] cpu_dout,

    input        cs,
    input [3:0]  cpu_addr,
    input cpu_rw,
    input [1:0] cpu_ds_n,

    input [13:0] color_in0 /* verilator public_flat */,
    input [13:0] color_in1 /* verilator public_flat */,
    input [13:0] color_in2 /* verilator public_flat */,
    output reg [13:0] color_out /* verilator public_flat */,

    ssbus_if.slave ssbus
);

reg [7:0] ctrl[16];

always_ff @(posedge clk) begin
    if (reset) begin
        int i;
        for (int i = 0; i < 16; i = i + 1) begin
            ctrl[i] <= 0;
        end
    end else begin
        if (cs) begin
            if (cpu_rw) begin
                cpu_dout <= { ctrl[cpu_addr[3:0]], ctrl[cpu_addr[3:0]] };
            end else begin
                if (~cpu_ds_n[0]) ctrl[cpu_addr[3:0]]  <= cpu_din[7:0];
            end
        end

        ssbus.setup(SS_IDX, 16, 0);
        if (ssbus.access(SS_IDX)) begin
            if (ssbus.write) begin
                ctrl[ssbus.addr[3:0]] <= ssbus.data[7:0];
                ssbus.write_ack(SS_IDX);
            end else if (ssbus.read) begin
                ssbus.read_response(SS_IDX, { 56'b0, ctrl[ssbus.addr[3:0]] });
            end
        end
    end
end


wire [1:0] sel0 = color_in0[13:12];
wire [1:0] sel1 = color_in1[13:12];
wire [1:0] sel2 = ctrl[1][7:6];

wire [15:0] prio_vals0 = { ctrl[5], ctrl[4] };
wire [15:0] prio_vals1 = { ctrl[7], ctrl[6] };
wire [15:0] prio_vals2 = { ctrl[9], ctrl[8] };

wire [3:0] prio0 = prio_vals0[ 4 * sel0 +: 4 ];
wire [3:0] prio1 = prio_vals1[ 4 * sel1 +: 4 ];
wire [3:0] prio2 = prio_vals2[ 4 * sel1 +: 4 ];

wire bm1 = ctrl[0][7] & ctrl[0][6]; 

always_ff @(posedge clk) begin
    if (ce_pixel) begin
        color_out <= color_in0;
        if (bm1 && (prio1 == (prio0 - 4'd1)) && |color_in1[3:0]) begin
            color_out <= { color_in1[13:4], color_in0[3:0] };
        end else if (bm1 && (prio1 == (prio0 + 4'd1)) && |color_in0[3:0]) begin
            color_out <= { color_in0[13:4], color_in1[3:0] };
        end else if (prio1 > prio0) begin
            if (prio2 > prio1) begin
                color_out <= color_in2;
            end else if (|color_in1[3:0]) begin
                color_out <= color_in1;
            end
        end else if (prio2 > prio0) begin
            color_out <= color_in2;
        end
    end
end


endmodule
